// Processor.v

// Generated using ACDS version 16.0 211

`timescale 1 ps / 1 ps
module Processor (
		input  wire       clk_clk,                   //      clk.clk
		output wire       done_writeresponsevalid_n, //     done.writeresponsevalid_n
		output wire [9:0] ledr_export,               //     ledr.export
		input  wire       reset_reset_n,             //    reset.reset_n
		input  wire       run_beginbursttransfer,    //      run.beginbursttransfer
		output wire [9:0] vgab_export,               //     vgab.export
		output wire       vgablank_export,           // vgablank.export
		output wire       vgaclk_export,             //   vgaclk.export
		output wire [9:0] vgag_export,               //     vgag.export
		output wire       vgahs_export,              //    vgahs.export
		output wire [9:0] vgar_export,               //     vgar.export
		output wire       vgasync_export,            //  vgasync.export
		output wire       vgavs_export               //    vgavs.export
	);

	wire  [31:0] processor_0_avalon_master_readdata;               // mm_interconnect_0:Processor_0_avalon_master_readdata -> Processor_0:DIN
	wire         processor_0_avalon_master_waitrequest;            // mm_interconnect_0:Processor_0_avalon_master_waitrequest -> Processor_0:waitrequest
	wire  [31:0] processor_0_avalon_master_address;                // Processor_0:Addr -> mm_interconnect_0:Processor_0_avalon_master_address
	wire   [3:0] processor_0_avalon_master_byteenable;             // Processor_0:byteenable -> mm_interconnect_0:Processor_0_avalon_master_byteenable
	wire         processor_0_avalon_master_read;                   // Processor_0:read -> mm_interconnect_0:Processor_0_avalon_master_read
	wire  [31:0] processor_0_avalon_master_writedata;              // Processor_0:DOUT -> mm_interconnect_0:Processor_0_avalon_master_writedata
	wire         processor_0_avalon_master_write;                  // Processor_0:write -> mm_interconnect_0:Processor_0_avalon_master_write
	wire         mm_interconnect_0_lda_0_s1_chipselect;            // mm_interconnect_0:LDA_0_s1_chipselect -> LDA_0:avs_s1_chipselect
	wire  [31:0] mm_interconnect_0_lda_0_s1_readdata;              // LDA_0:avs_s1_readdata -> mm_interconnect_0:LDA_0_s1_readdata
	wire         mm_interconnect_0_lda_0_s1_waitrequest;           // LDA_0:avs_s1_waitrequest -> mm_interconnect_0:LDA_0_s1_waitrequest
	wire   [2:0] mm_interconnect_0_lda_0_s1_address;               // mm_interconnect_0:LDA_0_s1_address -> LDA_0:avs_s1_address
	wire         mm_interconnect_0_lda_0_s1_read;                  // mm_interconnect_0:LDA_0_s1_read -> LDA_0:avs_s1_read
	wire         mm_interconnect_0_lda_0_s1_write;                 // mm_interconnect_0:LDA_0_s1_write -> LDA_0:avs_s1_write
	wire  [31:0] mm_interconnect_0_lda_0_s1_writedata;             // mm_interconnect_0:LDA_0_s1_writedata -> LDA_0:avs_s1_writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect; // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;   // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire   [7:0] mm_interconnect_0_onchip_memory2_0_s1_address;    // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable; // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;      // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;  // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;      // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         rst_controller_reset_out_reset;                   // rst_controller:reset_out -> [LDA_0:csi_clockreset_reset_n, Processor_0:reset, mm_interconnect_0:Processor_0_reset_reset_bridge_in_reset_reset, onchip_memory2_0:reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;               // rst_controller:reset_req -> [onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	wire y00;
	LDA_Peripheral lda_0 (
		.avs_s1_chipselect               (mm_interconnect_0_lda_0_s1_chipselect),  //               s1.chipselect
		.avs_s1_address                  (mm_interconnect_0_lda_0_s1_address),     //                 .address
		.avs_s1_read                     (mm_interconnect_0_lda_0_s1_read),        //                 .read
		.avs_s1_write                    (mm_interconnect_0_lda_0_s1_write),       //                 .write
		.avs_s1_writedata                (mm_interconnect_0_lda_0_s1_writedata),   //                 .writedata
		.avs_s1_readdata                 (mm_interconnect_0_lda_0_s1_readdata),    //                 .readdata
		.avs_s1_waitrequest              (mm_interconnect_0_lda_0_s1_waitrequest), //                 .waitrequest
		.coe_ledr_export_LEDR            (ledr_export),                            //             ledr.export
		.coe_vgar_export_VGA_R           (vgar_export),                            //             vgar.export
		.coe_vgag_export_VGA_G           (vgag_export),                            //             vgag.export
		.coe_vgab_export_VGA_B           (vgab_export),                            //             vgab.export
		.coe_vgahs_export_VGA_HS         (vgahs_export),                           //            vgahs.export
		.coe_vgavs_export_VGA_VS         (vgavs_export),                           //            vgavs.export
		.coe_vgablank_export_VGA_BLANK_N (vgablank_export),                        //         vgablank.export
		.coe_vgasync_export_VGA_SYNC_N   (vgasync_export),                         //          vgasync.export
		.coe_vgaclk_export_VGA_CLK       (vgaclk_export),                          //           vgaclk.export
		.csi_clockreset_clk              (clk_clk),                                //       clockreset.clk
		.csi_clockreset_reset_n          (~rst_controller_reset_out_reset),         // clockreset_reset.reset_n
		.y00 (y00)
	);

	wire [31:0] r1;
	proc processor_0 (
		.Addr        (processor_0_avalon_master_address),     // avalon_master.address
		.DIN         (processor_0_avalon_master_readdata),    //              .readdata
		.DOUT        (processor_0_avalon_master_writedata),   //              .writedata
		.byteenable  (processor_0_avalon_master_byteenable),  //              .byteenable
		.waitrequest (processor_0_avalon_master_waitrequest), //              .waitrequest
		.write       (processor_0_avalon_master_write),       //              .write
		.read        (processor_0_avalon_master_read),        //              .read
		.Clock       (clk_clk),                               //         clock.clk
		.Resetn       (~rst_controller_reset_out_reset),        //         reset.reset
		.Done        (done_writeresponsevalid_n),             //          Done.writeresponsevalid_n
		.Run         (run_beginbursttransfer),                 //           Run.beginbursttransfer
		.r1 (r1)
	);

	Processor_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)                //       .reset_req
	);

	Processor_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                 (clk_clk),                                          //                               clk_0_clk.clk
		.Processor_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                   // Processor_0_reset_reset_bridge_in_reset.reset
		.Processor_0_avalon_master_address             (processor_0_avalon_master_address),                //               Processor_0_avalon_master.address
		.Processor_0_avalon_master_waitrequest         (processor_0_avalon_master_waitrequest),            //                                        .waitrequest
		.Processor_0_avalon_master_byteenable          (processor_0_avalon_master_byteenable),             //                                        .byteenable
		.Processor_0_avalon_master_read                (processor_0_avalon_master_read),                   //                                        .read
		.Processor_0_avalon_master_readdata            (processor_0_avalon_master_readdata),               //                                        .readdata
		.Processor_0_avalon_master_write               (processor_0_avalon_master_write),                  //                                        .write
		.Processor_0_avalon_master_writedata           (processor_0_avalon_master_writedata),              //                                        .writedata
		.LDA_0_s1_address                              (mm_interconnect_0_lda_0_s1_address),               //                                LDA_0_s1.address
		.LDA_0_s1_write                                (mm_interconnect_0_lda_0_s1_write),                 //                                        .write
		.LDA_0_s1_read                                 (mm_interconnect_0_lda_0_s1_read),                  //                                        .read
		.LDA_0_s1_readdata                             (mm_interconnect_0_lda_0_s1_readdata),              //                                        .readdata
		.LDA_0_s1_writedata                            (mm_interconnect_0_lda_0_s1_writedata),             //                                        .writedata
		.LDA_0_s1_waitrequest                          (mm_interconnect_0_lda_0_s1_waitrequest),           //                                        .waitrequest
		.LDA_0_s1_chipselect                           (mm_interconnect_0_lda_0_s1_chipselect),            //                                        .chipselect
		.onchip_memory2_0_s1_address                   (mm_interconnect_0_onchip_memory2_0_s1_address),    //                     onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                     (mm_interconnect_0_onchip_memory2_0_s1_write),      //                                        .write
		.onchip_memory2_0_s1_readdata                  (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //                                        .readdata
		.onchip_memory2_0_s1_writedata                 (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //                                        .writedata
		.onchip_memory2_0_s1_byteenable                (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //                                        .byteenable
		.onchip_memory2_0_s1_chipselect                (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //                                        .chipselect
		.onchip_memory2_0_s1_clken                     (mm_interconnect_0_onchip_memory2_0_s1_clken)       //                                        .clken
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
